-- Code your testbench here
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

-- entity declaration for your testbench.Dont declare any ports here
ENTITY LPCMod_tb IS
END LPCMod_tb;

ARCHITECTURE behavior OF LPCMod_tb IS
   -- Component Declaration for the Unit Under Test (UUT)
    COMPONENT entity_lpcmod is  --'test' is the name of the module needed to be tested.
--just copy and paste the input and output ports of your module as such.
   port (
        pin_xbox_n_lrst     : in    std_logic;                      -- Xbox-side Reset signal
        pin_xbox_lclk       : in    std_logic;                      -- Xbox-side CLK, goes to flash chip too
        pin_pad_bt          : in    std_logic;                      -- Xbox power button. Labeled "BT" on silkscreen, near unrouted LCD pad array.
        pin_pad_h0          : in    std_logic;                      -- Unused pad? Labeled "H0" on silkscreen, near D0 pad. Will be used for flash bank switch (2 * 512KB).
        pout_flash_lframe   : out   std_logic;                      -- Only goes to flash chip. Is generated by code logic.
        pinout4_xbox_lad    : inout std_logic_vector(3 downto 0);   -- Xbox-side LPC IO
        pinout4_flash_lad   : inout std_logic_vector(3 downto 0);   -- Flash-side LPC IO
        pinout_pad_d0       : inout std_logic ;                     -- D0 control on Xbox motherbord. Useful on all motherboards but 1.6(b) should really USE L1 instead!
        pinout_pad_x        : inout std_logic;                      -- Supports D0 to sink in more current.
        pinout_pad_l1       : inout std_logic                       -- LFRAME control on the Motherboard. Useful only on 1.6(b)
    );
    END COMPONENT entity_lpcmod;
    
    signal pin_xbox_n_lrst : std_logic := '1';
    signal pin_xbox_lclk : std_logic := '0';
    signal pin_pad_bt : std_logic := '0';      --will stay 0 for this test.
    signal pin_pad_h0 : std_logic := 'Z';
    signal pout_flash_lframe : std_logic;
    signal pinout4_xbox_lad : std_logic_vector(3 downto 0) := "1111";
    signal pinout4_flash_lad : std_logic_vector(3 downto 0) := "0000";
    signal pinout_pad_d0 : std_logic := 'Z';
    signal pinout_pad_x  : std_logic := 'Z';
    signal pinout_pad_l1 : std_logic := 'Z';
    
    constant clk_period : time := 30 NS;
    
BEGIN
    -- Instantiate the Unit Under Test (UUT)
    uut: entity_lpcmod PORT MAP (
        pin_xbox_n_lrst,
        pin_xbox_lclk,
        pin_pad_bt,
        pin_pad_h0,
        pout_flash_lframe,
        pinout4_xbox_lad,
        pinout4_flash_lad,
        pinout_pad_d0,
        pinout_pad_x,
        pinout_pad_l1
    ); 
        
   -- Clock process definitions( clock with 50% duty cycle is generated here.
   clk_process :process
   begin
        pin_xbox_lclk <= '0';
        wait for clk_period/2;
        pin_xbox_lclk <= '1';
        wait for clk_period/2;
   end process;       
   
   
stim_proc: process
    begin    
        pin_xbox_n_lrst <= '0';
        pin_pad_bt <= '1';
        pinout_pad_d0 <= 'Z';
        pinout_pad_l1 <= 'Z';
        pin_pad_h0 <= '1';          --Flash write toggle. 0 for write disabled
        pinout4_flash_lad <= "ZZZZ";
        wait for clk_period;        --60 ns delay + 10 ns to shift new data entry. This make it so that new data is latched only 10ns before CLK rising edge.
        pin_pad_bt <= '0';         --Short PWR button press.
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        pin_pad_bt <= '1';
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        wait for 24 NS;         --Arbitrary delay induced on further data stimulation. In reality, the Xbox sets it's data for the next rising edge around 9 NS after the preceding rising edge of said data.
        pin_xbox_n_lrst <= '1';
        wait for clk_period;
        pin_pad_bt <= '0';
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --Start!
        wait for clk_period;
        pinout4_xbox_lad <= "0110"; --CYC
        wait for clk_period;
        pinout4_xbox_lad <= "1111"; --addr0
        wait for clk_period;
        pinout4_xbox_lad <= "1111"; --addr1
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --addr2
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --addr3
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr4
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr5
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr6
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr7
        wait for clk_period;
        pinout4_xbox_lad <= x"A";   --DATA1
        wait for clk_period;
        pinout4_xbox_lad <= x"A";   --DATA2
        wait for clk_period;
        pinout4_xbox_lad <= X"F";   --TARA1
        wait for clk_period;
        pinout4_xbox_lad <= "ZZZZ"; --TARA2
        pinout4_flash_lad <= X"F";
        wait for clk_period;
        pinout4_flash_lad <= "0000"; --SYNC
        wait for clk_period;
        pinout4_flash_lad <= X"F";   --TARB1
        wait for clk_period;
        pinout4_flash_lad <= "ZZZZ"; 
        pinout4_xbox_lad <= X"F";   --TARB2
        wait for clk_period;
        wait for clk_period;
        pin_pad_h0 <= '0';  -- Check that flash LFRAME isn't toggled on CYC Mem write ops
        wait for clk_period;
        wait for clk_period;
        
        
        
        pinout4_xbox_lad <= "0000"; --Start!
        wait for clk_period;
        pinout4_xbox_lad <= "0110"; --CYC
        wait for clk_period;
        pinout4_xbox_lad <= "1111"; --addr0
        wait for clk_period;
        pinout4_xbox_lad <= "1111"; --addr1
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --addr2
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --addr3
        wait for clk_period;
        pinout4_xbox_lad <= x"2";   --addr4
        wait for clk_period;
        pinout4_xbox_lad <= x"A";   --addr5
        wait for clk_period;
        pinout4_xbox_lad <= x"A";   --addr6
        wait for clk_period;
        pinout4_xbox_lad <= x"A";   --addr7
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --DATA1
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --DATA2
        wait for clk_period;
        pinout4_xbox_lad <= X"F";   --TARA1
        wait for clk_period;
        pinout4_xbox_lad <= "ZZZZ"; --TARA2
        pinout4_flash_lad <= X"F";
        wait for clk_period;
        pinout4_flash_lad <= "0000"; --SYNC
        wait for clk_period;
        pinout4_flash_lad <= X"F";   --TARB1
        wait for clk_period;
        pinout4_flash_lad <= "ZZZZ"; 
        pinout4_xbox_lad <= X"F";   --TARB2
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        
        
        
        pinout4_xbox_lad <= "0000"; --Start!
        wait for clk_period;
        pinout4_xbox_lad <= "0110"; --CYC
        wait for clk_period;
        pinout4_xbox_lad <= "1111"; --addr0
        wait for clk_period;
        pinout4_xbox_lad <= "1111"; --addr1
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --addr2
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --addr3
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr4
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr5
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr6
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr7
        wait for clk_period;
        pinout4_xbox_lad <= x"9";   --DATA1
        wait for clk_period;
        pinout4_xbox_lad <= x"0";   --DATA2
        wait for clk_period;
        pinout4_xbox_lad <= X"F";   --TARA1
        wait for clk_period;
        pinout4_xbox_lad <= "ZZZZ"; --TARA2
        pinout4_flash_lad <= X"F";
        wait for clk_period;
        pinout4_flash_lad <= "0000"; --SYNC
        wait for clk_period;
        pinout4_flash_lad <= X"F";   --TARB1
        wait for clk_period;
        pinout4_flash_lad <= "ZZZZ"; 
        pinout4_xbox_lad <= X"F";   --TARB2
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        
        
        
        pinout4_xbox_lad <= "0000"; --Start!
        wait for clk_period;
        pinout4_xbox_lad <= "0100"; --CYC
        wait for clk_period;
        pinout4_xbox_lad <= "1111"; --addr0
        wait for clk_period;
        pinout4_xbox_lad <= "1111"; --addr1
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --addr2
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --addr3
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr4
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr5
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr6
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr7
        wait for clk_period;
        pinout4_xbox_lad <= X"F";   --TARA1
        wait for clk_period;
        pinout4_xbox_lad <= "ZZZZ"; --TARA2
        pinout4_flash_lad <= X"F";
        wait for clk_period;
        pinout4_flash_lad <= "0000"; --SYNC
        wait for clk_period;
        pinout4_flash_lad <= x"2";   --DATA1
        wait for clk_period;
        pinout4_flash_lad <= x"5";   --DATA2
        wait for clk_period;
        pinout4_flash_lad <= X"F";   --TARB1
        wait for clk_period;
        pinout4_flash_lad <= "ZZZZ"; 
        pinout4_xbox_lad <= X"F";   --TARB2
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        
        
        
        pinout4_xbox_lad <= "0000"; --Start!
        wait for clk_period;
        pinout4_xbox_lad <= "0100"; --CYC
        wait for clk_period;
        pinout4_xbox_lad <= "1111"; --addr0
        wait for clk_period;
        pinout4_xbox_lad <= "1111"; --addr1
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --addr2
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --addr3
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr4
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr5
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr6
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr7
        wait for clk_period;
        pinout4_xbox_lad <= X"F";   --TARA1
        wait for clk_period;
        pinout4_xbox_lad <= "ZZZZ"; --TARA2
        pinout4_flash_lad <= X"F";
        wait for clk_period;
        pinout4_flash_lad <= "0000"; --SYNC
        wait for clk_period;
        pinout4_flash_lad <= x"F";   --DATA1
        wait for clk_period;
        pinout4_flash_lad <= x"B";   --DATA2
        wait for clk_period;
        pinout4_flash_lad <= X"F";   --TARB1
        wait for clk_period;
        pinout4_flash_lad <= "ZZZZ"; 
        pinout4_xbox_lad <= X"F";   --TARB2
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        
        
        
        pinout4_xbox_lad <= "0000"; --Start!
        wait for clk_period;
        pinout4_xbox_lad <= "0110"; --CYC
        wait for clk_period;
        pinout4_xbox_lad <= "1111"; --addr0
        wait for clk_period;
        pinout4_xbox_lad <= "1111"; --addr1
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --addr2
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --addr3
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr4
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr5
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr6
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr7
        wait for clk_period;
        pinout4_xbox_lad <= x"0";   --DATA1
        wait for clk_period;
        pinout4_xbox_lad <= x"F";   --DATA2
        wait for clk_period;
        pinout4_xbox_lad <= X"F";   --TARA1
        wait for clk_period;
        pinout4_xbox_lad <= "ZZZZ"; --TARA2
        pinout4_flash_lad <= X"F";
        wait for clk_period;
        pinout4_flash_lad <= "0000"; --SYNC
        wait for clk_period;
        pinout4_flash_lad <= X"F";   --TARB1
        wait for clk_period;
        pinout4_flash_lad <= "ZZZZ"; 
        pinout4_xbox_lad <= X"F";   --TARB2
        wait for clk_period;
        ASSERT FALSE REPORT "Test done." SEVERITY NOTE;
        wait;
    end process;

END behavior;
